`timescale 1ns / 1ps
module Imem(
		output [31:0] IW,
		input[15:0] pcOut);
	
	reg [31:0] M[0:65/*535*/];
	
	assign IW = M[pcOut];
	initial
	begin
		M[0] = 32'b10000000001010000000000000110010;
		M[1] = 32'b10000101011100000000000000000000;
		M[2] = 32'b00000000001010000000000001100100;
		M[3] = 32'b10101001101010000000000000000001;
		M[4] = 32'b10001001101110000000000000000001;
		M[5] = 32'b11010010000000000000000000010100;
		//M[26] = 32'b01010000001110000000000000000000;
		M[26] = 32'b00000000001110000000000001100100;
	end
endmodule
